msrss_no.v